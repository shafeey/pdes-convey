`define DW 32 	// Width of Event Data
`define TW 16		// Width of Timestamp
`define SIM_END_TIME 1000
